library verilog;
use verilog.vl_types.all;
entity inst_memory_vlg_vec_tst is
end inst_memory_vlg_vec_tst;
