library verilog;
use verilog.vl_types.all;
entity oac_lab2_vlg_vec_tst is
end oac_lab2_vlg_vec_tst;
